module SchoolSeatingSystem(input logic clk,
                           input logic [31:0] Student_No,
                           input logic [4:0] Seat_No,
                           input logic write,
                           output logic [10:0] time_out,
                           input logic [1:0] Seat_State);

   logic [10:0] setted_reset_time, setted_limit_time, Time;
   logic rst_temp;
   
   assign time_out = Time;
   
   set_up S0(setted_reset_time, setted_limit_time);
   TIMER T0(clk, setted_reset_time, rst_temp, Time);
   mem M0(rst_temp, write, Student_No, Time, Seat_State, Seat_No, setted_limit_time);
	
   
endmodule
