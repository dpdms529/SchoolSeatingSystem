module set_up(output logic [10:0] user_Reset_time,
         output logic [10:0] user_limit_time);
   assign user_Reset_time = 1440;
   assign user_limit_time = 10;
	
endmodule